module shift_rotate_2 (input CLK, SET, CLR, Sr_En, In, 
							output reg[3:0] q);
		


endmodule