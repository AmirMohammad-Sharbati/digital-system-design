module memory_tb ();


endmodule